module counter(
    
);
    
endmodule